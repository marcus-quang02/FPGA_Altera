
module PLL (
	clk_in_1_clk,
	reset_reset,
	clk_out_1_clk);	

	input		clk_in_1_clk;
	input		reset_reset;
	output		clk_out_1_clk;
endmodule
