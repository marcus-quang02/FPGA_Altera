
module pll (
	clk_50_clk,
	clk_out_clk,
	rst_reset);	

	input		clk_50_clk;
	output		clk_out_clk;
	input		rst_reset;
endmodule
